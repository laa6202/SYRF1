//phy_urx.v

module phy_urx(
uart_rx,
rx_data,
rx_vld,
//clk rst
clk_sys,
rst_n
);
output 				uart_rx;
input [31:0]	rx_data;
input 				rx_vld;
//clk rst
input clk_sys;
input rst_n;
//---------------------------------
//---------------------------------


endmodule
