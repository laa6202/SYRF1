//para_hit.v

module para_hit(
//data path
sm_data,
sm_vld,

//clk rst
clk_sys,
rst_n
);
//data path
input [15:0]	sm_data;
input					sm_vld;

input clk_sys;
input rst_n;
//--------------------------------
//--------------------------------



endmodule

