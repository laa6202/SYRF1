//fx_master.v

module fx_master(
tx_data,
tx_vld,
//clk rst
clk_sys,
rst_n
);
input [31:0]	tx_data;
input 				tx_vld;

//clk rst
input clk_sys;
input rst_n;
//--------------------------------------
//--------------------------------------



endmodule
