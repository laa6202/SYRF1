//fracture.v

module fracture(
//para input 
ph_ring,
ph_vld,
//register
cfg_ring_th,
stu_action,
clr_action,
//clk rst
clk_sys,
rst_n
);
//para input 
input [15:0]	ph_ring;
input					ph_vld;
//register
input [15:0]	cfg_ring_th;
output stu_action;
input  clr_action;
//clk rst
input clk_sys;
input rst_n;
//----------------------------------
//----------------------------------





endmodule

