//ad_filter.v

module ad_filter(
ad_data_s1,
ad_vld_s1,
ad_data_s2,
ad_vld_s2,
//clk rst
clk_sys,
rst_n
);
input [15:0]	ad_data_s1;
input					ad_vld_s1;
output [15:0]	ad_data_s2;
output				ad_vld_s2;
//clk rst
input	clk_sys;
input	rst_n;
//--------------------------------------
//--------------------------------------



endmodule

